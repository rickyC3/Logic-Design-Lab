`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/03/22 19:46:07
// Design Name: 
// Module Name: BCD_4bitsUpCnt
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module BCD_4bitsUpCnt(clk, rst, cnt);
input clk;
input rst;
output [11:0]cnt;
reg [3:0]inc;
endmodule
